library ieee;
use ieee.std_logic_1164.all;

entity controlador is
	Port(
		Resetn, clock: in std_logic;
		start, FinMem, Salir, Consultar_Saldo, Consultar_Mejores_Puntuaciones: in std_logic;
		HayTecla, CantValida, ApuestaValida, TermIntentos, t5s, NumValido, YaGano: in std_logic;
		esCaliente, esTibio, T2s, MayorMem, alcanzoN, Continuar: in std_logic;
		EnMem, LdMem, wr, EnInt, LdInt, En2s, Ld2s, En5s, Ld5s, EnVal: out std_logic;
		Ingrese, EnTecla, EnN, Sel, SelN, SelSumAP, EnSumAp, EnCant, Apuesta, EnAp, GetAlea, Adivine: out std_logic;
		EnMost, Caliente, Frio, Tibio, Perdio, Gano, SelSum, SelCant, EnDown, LdDown: out std_logic;
		SelAdd, SelMem, SelMost: out std_logic_vector(1 downto 0);
		est : out std_logic_vector(5 downTo 0);
		selNumber: out std_logic;
		Error: out std_logic
	);
end controlador;

Architecture sol of controlador is
	type estado is (T1, T2, T3, T4, T5, T6, T7, T8, T9, T10, T11, T12, T13, T14, T15, T16, T17, T18, T19, T20, T21, T22, T23, T24, T25, T26, T27, T28, T29, T30, T31, T32, T33, T34, T35, T36, T37,
						T38, T39, T40, T41, T42, T43, T44, T45, T46, T47, T48, T49, T50, T51,T52, T53, T54, T55, T56, T57, T58, T59, T60, T61, T62, T63, T64, t65, t66, t67, t68, t69);
	signal y: estado;

begin
-- Transiciones
Process(Resetn, clock)
Begin
	if Resetn = '0' then y <= T1;
	elsif clock'event and clock = '1' then
		case y is
			when T1 => y <= T2;
			when T2 => if FinMem = '0' then y<= T2; 
							else y<= T3; end if;
			when T3 => if start = '0' then y <= T3;
							else y<= T4; end if;
			when T4 => if start = '1' then y<= T4;
							else y<= T5; end if;
			when T5 => if Salir = '1' then y<= T3;
							elsif Consultar_Saldo = '1' then y<= T6;
							elsif Consultar_Mejores_Puntuaciones = '1' then y<= T7; 
							elsif HayTecla = '0' then y<= T5;
							else y<= T8; end if;
			when T6 => if Consultar_Saldo = '1' then y<= T6;
							else y<= T5; end if;
			when T7 => if Consultar_Mejores_Puntuaciones = '1' then y<= T7; else y <= T9; end if;
			when T8 => if HayTecla = '1' then y<= T8;
							else y<= T10; end if;
			when T9 => if T2s = '0' then y<= T9;
							elsif FinMem = '0' then y<= T9;
							else y <= T5; end if;
			when T10 => if salir = '1' then y<= T3;
							elsif Consultar_Saldo = '1' then y<= T11;
							elsif Consultar_Mejores_Puntuaciones = '1' then y<= T12; 
							elsif HayTecla = '0' then y<= T10;
							else y<= T13; end if;
			when T11 => if Consultar_Saldo = '1' then y<= T11;
							else y<= T10; end if;
			when T12 => if Consultar_Mejores_Puntuaciones = '1' then y<= T12; else y <= T14; end if;
			when T13 => if HayTecla = '1' then y<= T13;
							else y<= T15; end if;
			when T14 => if T2s = '0' then y<= T14; else y<= T64; end if;
			when T15 => y<= T16;
			when T16 => if salir = '1' then y<= T3;
							elsif Consultar_Saldo = '1' then y<= T17;
							elsif Consultar_Mejores_Puntuaciones = '1' then y<= T18; 
							elsif HayTecla = '0' then y<= T16;
							else y<= T19; end if;
			when T17 => if Consultar_Saldo = '1' then y<= T17;
							else y<= T16; end if;
			when T18 => if Consultar_Mejores_Puntuaciones = '1' then y<= T18; else y <= T20; end if;
			when T19 => if HayTecla = '1' then y<= T19;
							else y<=T21; end if;
			when T20 => if T2s = '0' then y<= T20;else y<= T65; end if;
			when T21 => y <= T22;
			when T22 => if cantValida = '0' then y<=T62;
							elsif continuar = '0' then y<= T22;
							else y<= T23; end if;
			when T23 => if salir = '1' then y<= T3;
							elsif Consultar_Saldo = '1' then y<= T24;
							elsif Consultar_Mejores_Puntuaciones = '1' then y<= T25; 
							elsif HayTecla = '0' then y<= T23;
							else y<= T26; end if;
			when T24 => if Consultar_Saldo = '1' then y<= T24;
							else y<= T23; end if;
			when T25 => if Consultar_Mejores_Puntuaciones = '1' then y<= T25; else y <= T27; end if;
			when T26 => if HayTecla = '1' then y<= T26;
							else y<=T28; end if;
			when T27 => if T2s = '0' then y<= T27; else y<= T66; end if;
			when T28 => if salir = '1' then y<= T3;
							elsif Consultar_Saldo = '1' then y<= T29;
							elsif Consultar_Mejores_Puntuaciones = '1' then y<= T30; 
							elsif HayTecla = '0' then y<= T28;
							else y<= T31; end if;
			when T29 => if Consultar_Saldo = '1' then y<= T29;
							else y<= T28; end if;
			when T30 => if Consultar_Mejores_Puntuaciones = '1' then y<= T30; else y <= T32; end if;
			when T31 => if HayTecla = '1' then y<= T31;
							else y<= T33; end if;
			when T32 => if T2s = '0' then y<= T32; else y<= T67; end if;
			when T33 => y<= T34;
			when T34 => if ApuestaValida = '0' then y<= T23;
							elsif Continuar = '0' then y<= T34;
							else y<= T35; end if;
			when T35 => y<= T36;
			when T36 => if TermIntentos = '1' then y<= T42;
							elsif salir = '1' then y<= T3;
							elsif Consultar_Saldo = '1' then y<= T37;
							elsif Consultar_Mejores_Puntuaciones = '1' then y<= T38; 
							elsif HayTecla = '0' then y<= T36;
							else y<= T39; end if;
			when T37 => if Consultar_Saldo = '1' then y<= T37;
							else y<= T36; end if;
			when T38 => if Consultar_Mejores_Puntuaciones = '1' then y<= T38; else y <= T40; end if;
			when T39 => if HayTecla = '1' then y<= T39;
							else y<= T41; end if;
			when T40 => if T2s = '0' then y<= T40; else y<= T68; end if;
			when T41 => if salir = '1' then y<= T3;
							elsif Consultar_Saldo = '1' then y<= T44;
							elsif Consultar_Mejores_Puntuaciones = '1' then y<= T45; 
							elsif HayTecla = '0' then y<= T41;
							else y<= T46; end if;
			when T42 => if T5s = '0' then y<= T42;
							else y<= T43; end if;
			when T43 => y<= T23;
			when T44 => if Consultar_Saldo = '1' then y<= T44;
							else y<= T41; end if;
			when T45 => if Consultar_Mejores_Puntuaciones = '1' then y<= T45; else y <= T47; end if;
			when T46 => if HayTecla = '1' then y<= T46;
							else y<= T48; end if;
			when T47 => if T2s = '0' then y<= T47; else y<= T69; end if;
			when T48 => y<= T49;
			when T49 => if NumValido = '0' then y<= T63;
							else y<= T50; end if;
			when T50 => if yaGano = '1' then y<= T51;
							elsif esCaliente = '1' then y<= T52;
							elsif esTibio = '1' then y<= T53;
							else y<= T54; end if;
			when T51 => if t5s = '0' then y<= T51;
							else y<= T55; end if;
			when T52 => if T2s = '0' then y<= T52;
							else y<= T36; end if;
			when T53 => if T2s = '0' then y<= T53;
							else y<= T36; end if;
			when T54 => if T2s = '0' then y<= T54;
							else y<= T36; end if;
			when T55 => y<= T56;
			when T56 => if FinMem = '1' then y<= T23;
							elsif MayorMem = '0' then y<= T56;
							else y<= T57; end if;
			when T57 => y<= T58;
			when T58 => y<= T59;
			when T59 => y<= T60;
			when T60 => if AlcanzoN = '0' then y<= T58;
							else y<= T61; end if;
			when T61=> y<= T23;
			when T62=> if T2s = '1' then y<= T5; end if;
			when T63=> if T2s = '1' then y<= T36; end if;
			when T64=> 	if FinMem = '0' then y<= T14;
							else y<= T10; end if;
			when T65=>  if FinMem = '0' then y<= T20;
							else y<= T16; end if;
			when T66=>  if FinMem = '0' then y<= T27;
							else y<= T23; end if;
			when T67=>  if FinMem = '0' then y<= T32;
							else y<= T28; end if;
			when T68=>  if FinMem = '0' then y<= T40;
							else y<= T36; end if;
			when T69=>  if FinMem = '0' then y<= T47;
							else y<= T41; end if;
		end case;
	end if;
end process;

--Salidas
Process(Resetn, clock, HayTecla, T5s, T2s)
begin
EnMem<='0'; LdMem<='0'; wr<='0'; EnInt<='0'; LdInt<='0'; SelSumAP<='0'; EnSumAp<= '0'; En2s<='0'; Ld2s<='0'; En5s<='0'; Ld5s<='0'; EnVal<='0';
EnMost<='0'; Caliente<='0'; Frio<='0'; Tibio<='0'; Perdio<='0'; Gano<='0'; SelSum<='0'; SelCant<='0'; EnDown<='0'; LdDown<='0';
Ingrese<='0'; EnTecla<='0'; EnN<='0'; Sel<='0'; SelN<='0'; EnCant<='0'; Apuesta<='0'; EnAp<='0'; GetAlea<='0'; Adivine<='0'; SelNumber <= '0'; Error <= '0';
SelAdd <= "00"; SelMem<= "00"; SelMost<= "00";
est <= "000000";
	case y is
		when T1 => Enmem <= '1'; LdMem<= '1'; EnTecla <= '1'; est <= "000001";
		when T2 => SelMem(0) <= '1'; EnMem <= '1'; Wr <= '1'; est <= "000010";
		when T3 => SelSumAP<='1'; EnSumAp<= '1'; EnInt<= '1'; LdInt<= '1'; En2s<= '1'; Ld2s<= '1'; En5s<= '1'; Ld5s<= '1'; EnN<='1';  est <= "000011";
		when T4 => est <= "000100";
		when T5 => Ingrese<= '1'; est <= "000101";
		when T6 => SelMost(1) <= '1'; EnMost<= '1'; est <= "000110";
		when T7 => EnMem <= '1'; LdMem <= '1'; est <= "000111";
		when T8 => if HayTecla ='1' then EnTecla<= '1'; EnN<= '1'; end if; est <= "001000";
		when T9 => En2s <= '1'; Ld2s <= '1'; EnMost <= '1'; SelMost(0)<= '1'; SelMost(1) <= '1'; est <= "001001";
						if(T2s = '1' and FinMem = '0') then EnMem <= '1'; end if;
		when T10 => Ingrese <= '1'; SelNumber <= '1'; EnMost <= '1'; est <= "001010";
		when T11 => SelMost(1) <= '1'; EnMost<= '1'; est <= "001011";
		when T12 => EnMem <= '1'; LdMem <= '1'; est <= "001100";
		when T13 => if HayTecla = '1' then EnTecla <= '1'; end if;est <= "001101";
		when T14 => En2s <= '1'; Ld2s <= '1'; EnMost <= '1'; SelMost(0)<= '1'; SelMost(1) <= '1'; est <= "001110";
		when T15 => EnN<= '1'; SelN<= '1'; est <= "001111";
		when T16 => Ingrese <= '1'; SelNumber <= '1'; EnMost <= '1'; est <= "010000";
		when T17 => SelMost(1) <= '1'; EnMost<= '1'; est <= "010001";
		when T18 => EnMem <= '1'; LdMem <= '1'; est <= "010010";
		when T19 => if HayTecla = '1' then EnTecla <= '1'; else EnN<= '1'; SelN<= '1'; end if; est <= "010011";
		when T20 => En2s <= '1'; Ld2s <= '1'; EnMost <= '1'; SelMost(0)<= '1'; SelMost(1) <= '1'; est <= "010100";
		when T21 => EnCant <= '1'; est <= "010101";
		when T22 => SelNumber <= '1'; EnMost <= '1'; est <= "010110";
		when T23 => Apuesta <= '1'; est <= "010111";
		when T24 => SelMost(1) <= '1'; EnMost<= '1'; est <= "011000";
		when T25 => EnMem <= '1'; LdMem <= '1'; est <= "011001";
		when T26 => if hayTecla = '1' then EnTecla <= '1'; EnN<= '1'; end if; est <= "011010";
		when T27 => En2s <= '1'; Ld2s <= '1'; EnMost <= '1'; SelMost(0)<= '1'; SelMost(1) <= '1'; est <= "011011";
		when T28 => Apuesta <= '1'; SelNumber <= '1'; EnMost <= '1'; est <= "011100";
		when T29 => SelMost(1) <= '1'; EnMost<= '1'; est <= "011101";
		when T30 => EnMem <= '1'; LdMem <= '1'; est <= "011110";
		when T31 => if HayTecla = '1' then EnTecla <= '1'; else EnN <= '1'; SelN <= '1'; end if; est <= "011111";
		when T32 => En2s <= '1'; Ld2s <= '1'; EnMost <= '1'; SelMost(0)<= '1'; SelMost(1) <= '1'; est <= "100000";						
		when T33 => EnAP <= '1'; est <= "100001";
		when T34 => EnMost <= '1'; selNumber <= '1'; est <= "100010";
		when T35 => GetAlea <= '1'; EnInt <= '1'; LdInt <= '1';est <= "100011";
		when T36 => Adivine <= '1'; EnMost <= '1';est <= "100100";
		when T37 => SelMost(1) <= '1'; EnMost<= '1'; est <= "100101";
		when T38 => EnMem <= '1'; LdMem <= '1'; est <= "100110";
		when T39 => EnMost <= '1';  est <= "100111";
						if HayTecla ='1' then EnTecla <= '1'; EnN <= '1'; end if;
		when T40 => En2s <= '1'; Ld2s <= '1'; EnMost <= '1'; SelMost(0)<= '1'; SelMost(1) <= '1'; est <= "101000";
		when T41 => Adivine <= '1'; EnMost <= '1'; est <= "101001";
		when T42 => Perdio <= '1'; EnMost <= '1'; En5s <= '1'; ld5s <= '1'; SelMost(0) <= '1'; est <= "101010";
						if t5s = '1' then En5s <= '1'; Ld5s <= '1'; end if;
		when T43 => SelSum <= '1'; SelCant <= '1'; EnCant <= '1'; est <= "101011";
		when T44 => SelMost(1) <= '1'; EnMost<= '1'; est <= "101100";
		when T45 => EnMem <= '1'; LdMem <= '1'; est <= "101101";
		when T46 => EnMost <= '1'; est <= "101110";
						if HayTecla = '1' then EnTecla <= '1'; end if;
		when T47 => En2s <= '1'; Ld2s <= '1'; EnMost <= '1'; SelMost(0)<= '1'; SelMost(1) <= '1'; est <= "101111";
		when T48 => EnN <= '1'; SelN <= '1'; est <= "110000";
		when T49 => EnMost <= '1'; est <= "110001";
		when T50 => EnMost <= '1'; est <= "110010";
		when T51 => Gano <= '1'; EnMost <= '1'; En5s <= '1'; ld5s <= '1'; SelMost(0) <= '1'; est <= "110011";
						if t5s = '1' then En5s <= '1'; ld5s <= '1'; end if;
		when T52 => Caliente <= '1'; En2s <= '1'; Ld2s <= '1'; est <= "110100";
						if T2s = '1' then En2s <= '1'; Ld2s <= '1'; EnInt <= '1'; end if;
		when T53 => Tibio <= '1'; En2s <= '1'; est <= "110101"; Ld2s <= '1';
						if T2s = '1' then En2s <= '1'; Ld2s <= '1'; EnInt <= '1'; end if;
		when T54 => Frio <= '1'; En2s <= '1'; est <= "110110"; Ld2s <= '1';
						if T2s = '1' then En2s <= '1'; Ld2s <= '1'; EnInt <= '1'; end if;
		when T55 => SelCant <= '1'; EnCant <= '1'; EnMem <= '1'; LdMem <= '1'; EnSumAp<='1'; est <= "110111";
		when T56 => EnMem <= '1'; est <= "111000";
		when T57 => EnDown <= '1'; LdDown <= '1';est <= "111001";
		when T58 => EnDown <= '1'; est <= "111010";
		when T59 => SelAdd(1) <= '1'; EnVal <= '1';est <= "111011";
		when T60 => SelAdd(0) <= '1'; SelMem(1) <= '1'; wr <= '1';est <= "111100";
		when T61 => wr <= '1'; est <= "111101";
		when T62 => Error <= '1'; En2s <= '1'; Ld2s <= '1'; if t2s = '1' then En2s <= '1'; Ld2s <= '1'; end if; est <= "111110";
		when T63 => Error <= '1'; En2s <= '1'; Ld2s <= '1'; if t2s = '1' then En2s <= '1'; Ld2s <= '1'; end if; est <= "111111";
		when T64 => EnMem <= '1';
		when T65 => EnMem <= '1';
		when T66 => EnMem <= '1';
		when T67 => EnMem <= '1';
		when T68 => EnMem <= '1';
		when T69 => EnMem <= '1';
	end case;
end process;

end sol;